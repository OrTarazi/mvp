
module HelloNios (
	clk_clk);	

	input		clk_clk;
endmodule
