// HelloNios.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module HelloNios (
		input  wire  clk_clk  // clk.clk
	);

	wire         hellonios_debug_reset_request_reset;                          // HelloNios:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] hellonios_data_master_readdata;                               // mm_interconnect_0:HelloNios_data_master_readdata -> HelloNios:d_readdata
	wire         hellonios_data_master_waitrequest;                            // mm_interconnect_0:HelloNios_data_master_waitrequest -> HelloNios:d_waitrequest
	wire         hellonios_data_master_debugaccess;                            // HelloNios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:HelloNios_data_master_debugaccess
	wire  [19:0] hellonios_data_master_address;                                // HelloNios:d_address -> mm_interconnect_0:HelloNios_data_master_address
	wire   [3:0] hellonios_data_master_byteenable;                             // HelloNios:d_byteenable -> mm_interconnect_0:HelloNios_data_master_byteenable
	wire         hellonios_data_master_read;                                   // HelloNios:d_read -> mm_interconnect_0:HelloNios_data_master_read
	wire         hellonios_data_master_write;                                  // HelloNios:d_write -> mm_interconnect_0:HelloNios_data_master_write
	wire  [31:0] hellonios_data_master_writedata;                              // HelloNios:d_writedata -> mm_interconnect_0:HelloNios_data_master_writedata
	wire  [31:0] hellonios_instruction_master_readdata;                        // mm_interconnect_0:HelloNios_instruction_master_readdata -> HelloNios:i_readdata
	wire         hellonios_instruction_master_waitrequest;                     // mm_interconnect_0:HelloNios_instruction_master_waitrequest -> HelloNios:i_waitrequest
	wire  [19:0] hellonios_instruction_master_address;                         // HelloNios:i_address -> mm_interconnect_0:HelloNios_instruction_master_address
	wire         hellonios_instruction_master_read;                            // HelloNios:i_read -> mm_interconnect_0:HelloNios_instruction_master_read
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;         // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;           // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest;        // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;            // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;               // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;              // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;          // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire  [31:0] mm_interconnect_0_mvp_accelerator_0_avalon_slave_0_readdata;  // mvp_accelerator_0:read_data -> mm_interconnect_0:mvp_accelerator_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_mvp_accelerator_0_avalon_slave_0_read;      // mm_interconnect_0:mvp_accelerator_0_avalon_slave_0_read -> mvp_accelerator_0:read
	wire         mm_interconnect_0_mvp_accelerator_0_avalon_slave_0_write;     // mm_interconnect_0:mvp_accelerator_0_avalon_slave_0_write -> mvp_accelerator_0:write
	wire  [31:0] mm_interconnect_0_mvp_accelerator_0_avalon_slave_0_writedata; // mm_interconnect_0:mvp_accelerator_0_avalon_slave_0_writedata -> mvp_accelerator_0:write_data
	wire  [31:0] mm_interconnect_0_hellonios_debug_mem_slave_readdata;         // HelloNios:debug_mem_slave_readdata -> mm_interconnect_0:HelloNios_debug_mem_slave_readdata
	wire         mm_interconnect_0_hellonios_debug_mem_slave_waitrequest;      // HelloNios:debug_mem_slave_waitrequest -> mm_interconnect_0:HelloNios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_hellonios_debug_mem_slave_debugaccess;      // mm_interconnect_0:HelloNios_debug_mem_slave_debugaccess -> HelloNios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_hellonios_debug_mem_slave_address;          // mm_interconnect_0:HelloNios_debug_mem_slave_address -> HelloNios:debug_mem_slave_address
	wire         mm_interconnect_0_hellonios_debug_mem_slave_read;             // mm_interconnect_0:HelloNios_debug_mem_slave_read -> HelloNios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_hellonios_debug_mem_slave_byteenable;       // mm_interconnect_0:HelloNios_debug_mem_slave_byteenable -> HelloNios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_hellonios_debug_mem_slave_write;            // mm_interconnect_0:HelloNios_debug_mem_slave_write -> HelloNios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_hellonios_debug_mem_slave_writedata;        // mm_interconnect_0:HelloNios_debug_mem_slave_writedata -> HelloNios:debug_mem_slave_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                         // mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                           // SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	wire  [15:0] mm_interconnect_0_sram_s1_address;                            // mm_interconnect_0:SRAM_s1_address -> SRAM:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                         // mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_s1_write;                              // mm_interconnect_0:SRAM_s1_write -> SRAM:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                          // mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	wire         mm_interconnect_0_sram_s1_clken;                              // mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                      // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                        // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [3:0] mm_interconnect_0_timer_0_s1_address;                         // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                           // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                       // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         irq_mapper_receiver0_irq;                                     // DEBUG:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] hellonios_irq_irq;                                            // irq_mapper:sender_irq -> HelloNios:irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [DEBUG:rst_n, HelloNios:reset_n, SRAM:reset, irq_mapper:reset, mm_interconnect_0:HelloNios_reset_reset_bridge_in_reset_reset, mvp_accelerator_0:resetn, rst_translator:in_reset, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [HelloNios:reset_req, SRAM:reset_req, rst_translator:reset_req_in]

	HelloNios_DEBUG debug (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                               //               irq.irq
	);

	HelloNios_HelloNios hellonios (
		.clk                                 (clk_clk),                                                 //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                         //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                      //                          .reset_req
		.d_address                           (hellonios_data_master_address),                           //               data_master.address
		.d_byteenable                        (hellonios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (hellonios_data_master_read),                              //                          .read
		.d_readdata                          (hellonios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (hellonios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (hellonios_data_master_write),                             //                          .write
		.d_writedata                         (hellonios_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (hellonios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (hellonios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (hellonios_instruction_master_read),                       //                          .read
		.i_readdata                          (hellonios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (hellonios_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (hellonios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (hellonios_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_hellonios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_hellonios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_hellonios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_hellonios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_hellonios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_hellonios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_hellonios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_hellonios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                         // custom_instruction_master.readra
	);

	HelloNios_SRAM sram (
		.clk        (clk_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                  // (terminated)
	);

	mvp_accelerator_avalon_slave mvp_accelerator_0 (
		.read       (mm_interconnect_0_mvp_accelerator_0_avalon_slave_0_read),      // avalon_slave_0.read
		.write      (mm_interconnect_0_mvp_accelerator_0_avalon_slave_0_write),     //               .write
		.write_data (mm_interconnect_0_mvp_accelerator_0_avalon_slave_0_writedata), //               .writedata
		.read_data  (mm_interconnect_0_mvp_accelerator_0_avalon_slave_0_readdata),  //               .readdata
		.clock      (clk_clk),                                                      //     clock_sink.clk
		.resetn     (~rst_controller_reset_out_reset)                               //     reset_sink.reset_n
	);

	HelloNios_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	HelloNios_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                               (clk_clk),                                                      //                             clk_0_clk.clk
		.HelloNios_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // HelloNios_reset_reset_bridge_in_reset.reset
		.HelloNios_data_master_address               (hellonios_data_master_address),                                //                 HelloNios_data_master.address
		.HelloNios_data_master_waitrequest           (hellonios_data_master_waitrequest),                            //                                      .waitrequest
		.HelloNios_data_master_byteenable            (hellonios_data_master_byteenable),                             //                                      .byteenable
		.HelloNios_data_master_read                  (hellonios_data_master_read),                                   //                                      .read
		.HelloNios_data_master_readdata              (hellonios_data_master_readdata),                               //                                      .readdata
		.HelloNios_data_master_write                 (hellonios_data_master_write),                                  //                                      .write
		.HelloNios_data_master_writedata             (hellonios_data_master_writedata),                              //                                      .writedata
		.HelloNios_data_master_debugaccess           (hellonios_data_master_debugaccess),                            //                                      .debugaccess
		.HelloNios_instruction_master_address        (hellonios_instruction_master_address),                         //          HelloNios_instruction_master.address
		.HelloNios_instruction_master_waitrequest    (hellonios_instruction_master_waitrequest),                     //                                      .waitrequest
		.HelloNios_instruction_master_read           (hellonios_instruction_master_read),                            //                                      .read
		.HelloNios_instruction_master_readdata       (hellonios_instruction_master_readdata),                        //                                      .readdata
		.DEBUG_avalon_jtag_slave_address             (mm_interconnect_0_debug_avalon_jtag_slave_address),            //               DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write               (mm_interconnect_0_debug_avalon_jtag_slave_write),              //                                      .write
		.DEBUG_avalon_jtag_slave_read                (mm_interconnect_0_debug_avalon_jtag_slave_read),               //                                      .read
		.DEBUG_avalon_jtag_slave_readdata            (mm_interconnect_0_debug_avalon_jtag_slave_readdata),           //                                      .readdata
		.DEBUG_avalon_jtag_slave_writedata           (mm_interconnect_0_debug_avalon_jtag_slave_writedata),          //                                      .writedata
		.DEBUG_avalon_jtag_slave_waitrequest         (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest),        //                                      .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect          (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),         //                                      .chipselect
		.HelloNios_debug_mem_slave_address           (mm_interconnect_0_hellonios_debug_mem_slave_address),          //             HelloNios_debug_mem_slave.address
		.HelloNios_debug_mem_slave_write             (mm_interconnect_0_hellonios_debug_mem_slave_write),            //                                      .write
		.HelloNios_debug_mem_slave_read              (mm_interconnect_0_hellonios_debug_mem_slave_read),             //                                      .read
		.HelloNios_debug_mem_slave_readdata          (mm_interconnect_0_hellonios_debug_mem_slave_readdata),         //                                      .readdata
		.HelloNios_debug_mem_slave_writedata         (mm_interconnect_0_hellonios_debug_mem_slave_writedata),        //                                      .writedata
		.HelloNios_debug_mem_slave_byteenable        (mm_interconnect_0_hellonios_debug_mem_slave_byteenable),       //                                      .byteenable
		.HelloNios_debug_mem_slave_waitrequest       (mm_interconnect_0_hellonios_debug_mem_slave_waitrequest),      //                                      .waitrequest
		.HelloNios_debug_mem_slave_debugaccess       (mm_interconnect_0_hellonios_debug_mem_slave_debugaccess),      //                                      .debugaccess
		.mvp_accelerator_0_avalon_slave_0_write      (mm_interconnect_0_mvp_accelerator_0_avalon_slave_0_write),     //      mvp_accelerator_0_avalon_slave_0.write
		.mvp_accelerator_0_avalon_slave_0_read       (mm_interconnect_0_mvp_accelerator_0_avalon_slave_0_read),      //                                      .read
		.mvp_accelerator_0_avalon_slave_0_readdata   (mm_interconnect_0_mvp_accelerator_0_avalon_slave_0_readdata),  //                                      .readdata
		.mvp_accelerator_0_avalon_slave_0_writedata  (mm_interconnect_0_mvp_accelerator_0_avalon_slave_0_writedata), //                                      .writedata
		.SRAM_s1_address                             (mm_interconnect_0_sram_s1_address),                            //                               SRAM_s1.address
		.SRAM_s1_write                               (mm_interconnect_0_sram_s1_write),                              //                                      .write
		.SRAM_s1_readdata                            (mm_interconnect_0_sram_s1_readdata),                           //                                      .readdata
		.SRAM_s1_writedata                           (mm_interconnect_0_sram_s1_writedata),                          //                                      .writedata
		.SRAM_s1_byteenable                          (mm_interconnect_0_sram_s1_byteenable),                         //                                      .byteenable
		.SRAM_s1_chipselect                          (mm_interconnect_0_sram_s1_chipselect),                         //                                      .chipselect
		.SRAM_s1_clken                               (mm_interconnect_0_sram_s1_clken),                              //                                      .clken
		.timer_0_s1_address                          (mm_interconnect_0_timer_0_s1_address),                         //                            timer_0_s1.address
		.timer_0_s1_write                            (mm_interconnect_0_timer_0_s1_write),                           //                                      .write
		.timer_0_s1_readdata                         (mm_interconnect_0_timer_0_s1_readdata),                        //                                      .readdata
		.timer_0_s1_writedata                        (mm_interconnect_0_timer_0_s1_writedata),                       //                                      .writedata
		.timer_0_s1_chipselect                       (mm_interconnect_0_timer_0_s1_chipselect)                       //                                      .chipselect
	);

	HelloNios_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (hellonios_irq_irq)               //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (hellonios_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_in1      (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
